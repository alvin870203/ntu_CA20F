module MUX# (
    parameter DATA_WIDTH = 32
)(
    
);